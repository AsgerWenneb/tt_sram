magic
tech sky130B
magscale 1 2
timestamp 1740166019
<< nwell >>
rect 22728 21744 23050 22052
<< nmos >>
rect 22858 21446 22918 21538
<< pmos >>
rect 22858 21780 22918 21870
<< ndiff >>
rect 22768 21528 22858 21538
rect 22768 21474 22784 21528
rect 22838 21474 22858 21528
rect 22768 21446 22858 21474
rect 22918 21524 23006 21538
rect 22918 21472 22932 21524
rect 22984 21472 23006 21524
rect 22918 21446 23006 21472
<< pdiff >>
rect 22764 21856 22858 21870
rect 22764 21798 22782 21856
rect 22832 21798 22858 21856
rect 22764 21780 22858 21798
rect 22918 21858 23014 21870
rect 22918 21792 22932 21858
rect 22996 21792 23014 21858
rect 22918 21780 23014 21792
<< ndiffc >>
rect 22784 21474 22838 21528
rect 22932 21472 22984 21524
<< pdiffc >>
rect 22782 21798 22832 21856
rect 22932 21792 22996 21858
<< psubdiff >>
rect 22812 21234 22836 21296
rect 22908 21234 22932 21296
<< nsubdiff >>
rect 22776 21942 22800 22004
rect 22868 21942 22892 22004
<< psubdiffcont >>
rect 22836 21234 22908 21296
<< nsubdiffcont >>
rect 22800 21942 22868 22004
<< poly >>
rect 22858 21870 22918 21900
rect 22858 21720 22918 21780
rect 22738 21700 22918 21720
rect 22738 21626 22764 21700
rect 22836 21626 22918 21700
rect 22738 21600 22918 21626
rect 22858 21538 22918 21600
rect 22858 21420 22918 21446
<< polycont >>
rect 22764 21626 22836 21700
<< locali >>
rect 22560 22004 23048 22042
rect 22560 21948 22588 22004
rect 22666 21948 22800 22004
rect 22560 21942 22800 21948
rect 22868 21942 23048 22004
rect 22560 21912 23048 21942
rect 22560 21910 22834 21912
rect 22782 21856 22834 21910
rect 22932 21858 22996 21874
rect 22782 21782 22832 21798
rect 22932 21776 22996 21792
rect 22748 21626 22764 21700
rect 22836 21626 22854 21700
rect 22932 21676 22984 21776
rect 22932 21632 22942 21676
rect 22976 21632 22984 21676
rect 22784 21528 22838 21546
rect 22784 21458 22838 21474
rect 22932 21524 22984 21632
rect 22784 21340 22836 21458
rect 22932 21456 22984 21472
rect 22616 21298 23108 21340
rect 22616 21230 22658 21298
rect 22742 21296 23108 21298
rect 22742 21234 22836 21296
rect 22908 21234 23108 21296
rect 22742 21230 23108 21234
rect 22616 21196 23108 21230
<< viali >>
rect 22588 21948 22666 22004
rect 22780 21644 22820 21684
rect 22942 21632 22976 21676
rect 22658 21230 22742 21298
<< metal1 >>
rect 22450 22004 22696 22030
rect 22450 21948 22588 22004
rect 22666 21948 22696 22004
rect 204 21882 534 21936
rect 22450 21924 22696 21948
rect 204 21702 250 21882
rect 490 21878 534 21882
rect 490 21876 18230 21878
rect 22452 21876 22542 21924
rect 490 21748 22542 21876
rect 490 21702 18230 21748
rect 204 21670 18230 21702
rect 22762 21696 22838 21702
rect 204 21662 534 21670
rect 18816 21662 18884 21666
rect 18816 21610 18826 21662
rect 18878 21659 18884 21662
rect 22762 21659 22768 21696
rect 18878 21632 22768 21659
rect 22832 21659 22838 21696
rect 22928 21676 22990 21690
rect 22928 21659 22942 21676
rect 22832 21632 22942 21659
rect 22976 21659 22990 21676
rect 22976 21632 23039 21659
rect 18878 21631 23039 21632
rect 18878 21610 18884 21631
rect 22762 21626 22838 21631
rect 22928 21618 22990 21631
rect 18816 21602 18884 21610
rect 22630 21318 22782 21326
rect 900 21298 22782 21318
rect 900 21292 22658 21298
rect 900 21228 932 21292
rect 1006 21230 22658 21292
rect 22742 21230 22782 21298
rect 1006 21228 22782 21230
rect 900 21198 22782 21228
<< via1 >>
rect 250 21702 490 21882
rect 18826 21610 18878 21662
rect 22768 21684 22832 21696
rect 22768 21644 22780 21684
rect 22780 21644 22820 21684
rect 22820 21644 22832 21684
rect 22768 21632 22832 21644
rect 932 21228 1006 21292
<< metal2 >>
rect 204 21890 540 21936
rect 204 21882 256 21890
rect 476 21882 540 21890
rect 204 21702 250 21882
rect 490 21702 540 21882
rect 204 21660 540 21702
rect 22758 21696 22844 21706
rect 18806 21662 18898 21676
rect 18806 21604 18826 21662
rect 18878 21660 18898 21662
rect 18882 21604 18898 21660
rect 22758 21632 22768 21696
rect 22832 21632 22844 21696
rect 22758 21622 22844 21632
rect 18806 21588 18898 21604
rect 860 21300 1068 21346
rect 860 21202 912 21300
rect 1010 21202 1068 21300
rect 860 21162 1068 21202
<< via2 >>
rect 256 21882 476 21890
rect 256 21724 476 21882
rect 18826 21610 18878 21660
rect 18878 21610 18882 21660
rect 18826 21604 18882 21610
rect 22768 21632 22832 21696
rect 912 21292 1010 21300
rect 912 21228 932 21292
rect 932 21228 1006 21292
rect 1006 21228 1010 21292
rect 912 21202 1010 21228
<< metal3 >>
rect 23812 22020 23890 22026
rect 23812 21956 23818 22020
rect 23884 21956 23890 22020
rect 198 21922 544 21954
rect 23812 21948 23890 21956
rect 198 21708 252 21922
rect 492 21708 544 21922
rect 198 21664 544 21708
rect 22742 21696 22858 21720
rect 18790 21678 18924 21696
rect 18790 21586 18808 21678
rect 18904 21586 18924 21678
rect 22742 21663 22768 21696
rect 18790 21570 18924 21586
rect 22380 21632 22768 21663
rect 22832 21632 22858 21696
rect 22380 21603 22858 21632
rect 858 21310 1068 21350
rect 858 21204 898 21310
rect 1012 21204 1068 21310
rect 858 21202 912 21204
rect 1010 21202 1068 21204
rect 858 21158 1068 21202
rect 22380 21062 22440 21603
rect 22742 21602 22858 21603
rect 23818 21062 23878 21948
rect 22380 21002 23878 21062
<< via3 >>
rect 23818 21956 23884 22020
rect 252 21890 492 21922
rect 252 21724 256 21890
rect 256 21724 476 21890
rect 476 21724 492 21890
rect 252 21708 492 21724
rect 18808 21660 18904 21678
rect 18808 21604 18826 21660
rect 18826 21604 18882 21660
rect 18882 21604 18904 21660
rect 18808 21586 18904 21604
rect 898 21300 1012 21310
rect 898 21204 912 21300
rect 912 21204 1010 21300
rect 1010 21204 1012 21300
<< metal4 >>
rect 6134 22104 6194 22304
rect 6686 22104 6746 22304
rect 7238 22104 7298 22304
rect 7790 22104 7850 22304
rect 8342 22104 8402 22304
rect 8894 22104 8954 22304
rect 9446 22104 9506 22304
rect 9998 22104 10058 22304
rect 10550 22104 10610 22304
rect 11102 22104 11162 22304
rect 11654 22104 11714 22304
rect 12206 22104 12266 22304
rect 12758 22104 12818 22304
rect 13310 22104 13370 22304
rect 13862 22104 13922 22304
rect 14414 22104 14474 22304
rect 14966 22104 15026 22304
rect 15518 22104 15578 22304
rect 16070 22104 16130 22304
rect 16622 22104 16682 22304
rect 17174 22104 17234 22304
rect 17726 22104 17786 22304
rect 18278 22104 18338 22304
rect 200 21922 600 22000
rect 200 21708 252 21922
rect 492 21708 600 21922
rect 200 1000 600 21708
rect 800 21310 1200 22000
rect 18830 21696 18890 22304
rect 19382 22104 19442 22304
rect 19934 22104 19994 22304
rect 20486 22104 20546 22304
rect 21038 22104 21098 22304
rect 21590 22104 21650 22304
rect 22142 22104 22202 22304
rect 22694 22104 22754 22304
rect 23246 21724 23306 22304
rect 23798 22032 23858 22304
rect 24350 22104 24410 22304
rect 24902 22104 24962 22304
rect 25454 22104 25514 22304
rect 26006 22104 26066 22304
rect 26558 22104 26618 22304
rect 27110 22104 27170 22304
rect 27662 22104 27722 22304
rect 28214 22104 28274 22304
rect 28766 22104 28826 22304
rect 29318 22104 29378 22304
rect 23798 22020 23900 22032
rect 23798 21956 23818 22020
rect 23884 21956 23900 22020
rect 23798 21942 23900 21956
rect 18790 21678 18920 21696
rect 18790 21586 18808 21678
rect 18904 21586 18920 21678
rect 18790 21572 18920 21586
rect 800 21204 898 21310
rect 1012 21204 1200 21310
rect 800 1000 1200 21204
<< labels >>
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 22104 29378 22304 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 22104 28274 22304 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27662 22104 27722 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 27110 22104 27170 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 26006 22104 26066 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 25454 22104 25514 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 24902 22104 24962 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 23798 22104 23858 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 23246 22104 23306 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 22694 22104 22754 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 21590 22104 21650 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 21038 22104 21098 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 20486 22104 20546 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19382 22104 19442 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 9998 22104 10058 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal output
flabel metal4 s 9446 22104 9506 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal output
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal output
flabel metal4 s 8342 22104 8402 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal output
flabel metal4 s 7790 22104 7850 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal output
flabel metal4 s 7238 22104 7298 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal output
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal output
flabel metal4 s 6134 22104 6194 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal output
flabel metal4 s 14414 22104 14474 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal output
flabel metal4 s 13862 22104 13922 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal output
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal output
flabel metal4 s 12758 22104 12818 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal output
flabel metal4 s 12206 22104 12266 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal output
flabel metal4 s 11654 22104 11714 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal output
flabel metal4 s 10550 22104 10610 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal output
flabel metal4 s 18830 22104 18890 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal output
flabel metal4 s 18278 22104 18338 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal output
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal output
flabel metal4 s 17174 22104 17234 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal output
flabel metal4 s 16622 22104 16682 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal output
flabel metal4 s 16070 22104 16130 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal output
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal output
flabel metal4 s 14966 22104 15026 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal output
flabel metal4 200 1000 600 22000 1 FreeSans 400 0 0 0 VDPWR
port 43 nsew power bidirectional
flabel metal4 800 1000 1200 22000 1 FreeSans 400 0 0 0 VGND
port 44 nsew ground bidirectional
rlabel polycont 22800 21664 22800 21664 1 A
rlabel viali 22958 21666 22958 21666 1 Y
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
