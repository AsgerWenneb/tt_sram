magic
tech sky130A
magscale 1 2
timestamp 1741791709
<< nwell >>
rect -189 94 110 262
<< nmos >>
rect -15 -73 15 11
<< pmos >>
rect -15 130 15 214
<< ndiff >>
rect -75 -1 -15 11
rect -75 -61 -61 -1
rect -27 -61 -15 -1
rect -75 -73 -15 -61
rect 15 -1 73 11
rect 15 -61 27 -1
rect 61 -61 73 -1
rect 15 -73 73 -61
<< pdiff >>
rect -75 202 -15 214
rect -75 142 -61 202
rect -27 142 -15 202
rect -75 130 -15 142
rect 15 202 73 214
rect 15 142 27 202
rect 61 142 73 202
rect 15 130 73 142
<< ndiffc >>
rect -61 -61 -27 -1
rect 27 -61 61 -1
<< pdiffc >>
rect -61 142 -27 202
rect 27 142 61 202
<< psubdiff >>
rect -153 -1 -75 11
rect -153 -61 -129 -1
rect -95 -61 -75 -1
rect -153 -73 -75 -61
<< nsubdiff >>
rect -153 202 -75 214
rect -153 142 -129 202
rect -95 142 -75 202
rect -153 130 -75 142
<< psubdiffcont >>
rect -129 -61 -95 -1
<< nsubdiffcont >>
rect -129 142 -95 202
<< poly >>
rect -15 214 15 240
rect -15 99 15 130
rect -33 83 33 99
rect -33 49 -17 83
rect 17 49 33 83
rect -33 33 33 49
rect -15 11 15 33
rect -15 -99 15 -73
<< polycont >>
rect -17 49 17 83
<< locali >>
rect -129 202 -27 218
rect -95 142 -61 202
rect -129 126 -27 142
rect 27 202 61 218
rect 61 142 110 160
rect 27 126 110 142
rect -189 49 -17 83
rect 17 49 33 83
rect 76 15 110 126
rect -129 -1 -27 15
rect -95 -61 -61 -1
rect -129 -77 -27 -61
rect 27 -1 110 15
rect 61 -19 110 -1
rect 27 -77 61 -61
<< viali >>
rect -129 142 -95 202
<< metal1 >>
rect -189 202 -89 214
rect -189 142 -129 202
rect -95 142 -89 202
rect -189 130 -89 142
rect -189 -73 -89 11
<< labels >>
rlabel locali -189 66 -189 66 7 A
port 1 w
rlabel locali 110 66 110 66 3 X
port 2 e
rlabel metal1 -189 -31 -189 -31 7 VGND
port 3 w
rlabel metal1 -189 172 -189 172 7 VPWR
port 4 w
<< properties >>
string FIXED_BBOX 0 0 100 100
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
