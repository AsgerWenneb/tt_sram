MACRO my_inverter
  CLASS BLOCK ;
  FOREIGN my_inverter ;
  ORIGIN 0.945 0.495 ;
  SIZE 1.495 BY 1.805 ;
  PIN A
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT -0.945 0.245 0.165 0.415 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA 0.243600 ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.800 0.305 1.090 ;
        RECT 0.135 0.630 0.550 0.800 ;
        RECT 0.380 0.075 0.550 0.630 ;
        RECT 0.135 -0.095 0.550 0.075 ;
        RECT 0.135 -0.385 0.305 -0.095 ;
    END
  END X
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.945 -0.365 -0.445 0.055 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT -0.945 0.650 -0.445 1.070 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT -0.645 -0.385 -0.135 0.075 ;
  END
END my_inverter
END LIBRARY

