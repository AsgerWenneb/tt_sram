magic
tech sky130A
magscale 1 2
timestamp 1741186866
<< nwell >>
rect -180 150 150 340
<< nmos >>
rect 10 -60 40 30
<< pmos >>
rect 10 200 40 290
<< ndiff >>
rect -60 10 10 30
rect -60 -40 -40 10
rect -6 -40 10 10
rect -60 -60 10 -40
rect 40 10 110 30
rect 40 -40 60 10
rect 94 -40 110 10
rect 40 -60 110 -40
<< pdiff >>
rect -60 270 10 290
rect -60 220 -40 270
rect -6 220 10 270
rect -60 200 10 220
rect 40 270 110 290
rect 40 220 60 270
rect 100 220 110 270
rect 40 200 110 220
<< ndiffc >>
rect -40 -40 -6 10
rect 60 -40 94 10
<< pdiffc >>
rect -40 220 -6 270
rect 60 220 100 270
<< psubdiff >>
rect -140 30 -85 40
rect -140 10 -60 30
rect -140 -40 -110 10
rect -76 -40 -60 10
rect -140 -60 -60 -40
rect -140 -70 -85 -60
<< nsubdiff >>
rect -140 290 -85 300
rect -140 270 -60 290
rect -140 220 -120 270
rect -80 220 -60 270
rect -140 200 -60 220
rect -140 190 -85 200
<< psubdiffcont >>
rect -110 -40 -76 10
<< nsubdiffcont >>
rect -120 220 -80 270
<< poly >>
rect 10 290 40 320
rect -110 124 -40 140
rect -110 90 -90 124
rect -56 120 -40 124
rect 10 120 40 200
rect -56 90 40 120
rect -110 70 -40 90
rect 10 30 40 90
rect 10 -86 40 -60
<< polycont >>
rect -90 90 -56 124
<< locali >>
rect -180 270 10 290
rect -180 220 -120 270
rect -80 220 -40 270
rect -6 220 10 270
rect -180 200 10 220
rect 50 270 110 290
rect 50 220 60 270
rect 100 220 110 270
rect 50 140 110 220
rect -180 124 -40 140
rect -180 90 -90 124
rect -56 90 -40 124
rect -180 70 -40 90
rect 50 70 150 140
rect -180 10 10 30
rect -180 -40 -110 10
rect -76 -40 -40 10
rect -6 -40 10 10
rect -180 -60 10 -40
rect 50 10 110 70
rect 50 -40 60 10
rect 94 -40 110 10
rect 50 -60 110 -40
<< labels >>
rlabel locali -180 110 -180 110 7 A
port 1 w
rlabel locali -180 250 -180 250 7 VP
port 2 w
rlabel locali -180 -10 -180 -10 7 VN
port 3 w
rlabel locali 150 110 150 110 3 Y
port 4 e
<< end >>
