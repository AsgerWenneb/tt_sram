VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO invering_buffer
  CLASS BLOCK ;
  FOREIGN invering_buffer ;
  ORIGIN 0.800 0.150 ;
  SIZE 1.200 BY 1.000 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT -0.945 0.245 0.165 0.415 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.243600 ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.800 0.305 1.090 ;
        RECT 0.135 0.630 0.550 0.800 ;
        RECT 0.380 0.075 0.550 0.630 ;
        RECT 0.135 -0.095 0.550 0.075 ;
        RECT 0.135 -0.385 0.305 -0.095 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.945 -0.365 -0.445 0.055 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.945 0.470 0.550 1.310 ;
      LAYER li1 ;
        RECT -0.645 0.630 -0.135 1.090 ;
      LAYER met1 ;
        RECT -0.945 0.650 -0.445 1.070 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT -0.645 -0.385 -0.135 0.075 ;
  END
END invering_buffer
END LIBRARY

